library verilog;
use verilog.vl_types.all;
entity alu32Testbench is
end alu32Testbench;
