library verilog;
use verilog.vl_types.all;
entity andTestbench is
end andTestbench;
