module mult32(input [31:0]multiplier, multiplicand, output product);

/*
wire[2:0] s,n;
wire go ,is_less ,write, add, sr;

initial begin
product[31:0] =  multiplier;
end

controller(s, product[0],go,is_less, add, sr,write, n);

always @(*)begin
	if(sr)begin
		product <= (product >> 1);
	end
end	
*/
endmodule
