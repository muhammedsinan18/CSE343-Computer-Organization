library verilog;
use verilog.vl_types.all;
entity sltTestbench is
end sltTestbench;
