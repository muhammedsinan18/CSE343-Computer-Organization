library verilog;
use verilog.vl_types.all;
entity xorTestbench is
end xorTestbench;
