library verilog;
use verilog.vl_types.all;
entity orTestbench is
end orTestbench;
