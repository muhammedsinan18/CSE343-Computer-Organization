library verilog;
use verilog.vl_types.all;
entity addTestbench is
end addTestbench;
