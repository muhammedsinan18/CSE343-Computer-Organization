library verilog;
use verilog.vl_types.all;
entity subTestbench is
end subTestbench;
