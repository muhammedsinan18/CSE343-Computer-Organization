library verilog;
use verilog.vl_types.all;
entity norTestbench is
end norTestbench;
